module Multiplier(
    input signed [31:0] A, B,
    output signed [63:0] P
);

    // TODO: implement Multiplier here
    // Note: Do NOT use built-in operator * here.
    always @(*) begin
        // TODO
    end

endmodule
